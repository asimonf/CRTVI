package Utils is
   type PixelParam is (M, N, C, K);
end package Utils;